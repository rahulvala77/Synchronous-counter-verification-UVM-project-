//-------------------------------------------------------
//file-name -> counter_parameters.sv
//class -> NA 
//methods ->  NA
//description -> parameters declaraed in this file 
//-------------------------------------------------------
parameter n = 2;

parameter number =2;

parameter int unsigned RESET_MIN=19;
parameter int unsigned RESET_MAX=20; 
